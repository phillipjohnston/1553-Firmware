----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    20:33:34 11/07/2012 
-- Design Name: 
-- Module Name:    SIGNAL_PLACEHOLDER - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity SIGNAL_PLACEHOLDER is
	PORT(
		EXP_IO_0 : OUT STD_LOGIC;
		EXP_IO_1 : OUT STD_LOGIC;
		EXP_IO_2 : OUT STD_LOGIC;
		EXP_IO_3 : OUT STD_LOGIC;
		EXP_IO_4 : OUT STD_LOGIC;
		EXP_IO_5 : OUT STD_LOGIC;
		EXP_IO_6 : OUT STD_LOGIC;
		EXP_IO_7 : OUT STD_LOGIC;
		EXP_IO_8 : OUT STD_LOGIC;
		EXP_IO_9 : OUT STD_LOGIC;
		EXP_IO_10 : OUT STD_LOGIC;
		EXP_IO_11 : OUT STD_LOGIC;
		EXP_IO_12 : OUT STD_LOGIC;
		EXP_IO_13 : OUT STD_LOGIC;
		
		MTRUN : OUT STD_LOGIC;
		RT1ENA : OUT STD_LOGIC;
		BCTRIG : OUT STD_LOGIC;
		TXINHB : OUT STD_LOGIC;
		TXINHA : OUT STD_LOGIC;
		ACTIVE : OUT STD_LOGIC;
		READY : OUT STD_LOGIC;
		ACKIRQ : OUT STD_LOGIC;
		nIRQ : OUT STD_LOGIC;
		nRT1MC8 : OUT STD_LOGIC;
		MTPKRDY : OUT STD_LOGIC;
		RT1SSF : OUT STD_LOGIC;
		BCENA : OUT STD_LOGIC;
		TEST : OUT STD_LOGIC;
		
		
		
	);
end SIGNAL_PLACEHOLDER;

architecture Behavioral of SIGNAL_PLACEHOLDER is

begin


end Behavioral;

